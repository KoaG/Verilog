module mux4to1_bh_tb();

reg [3:0]i;
reg [1:0]sel;
wire y;

mux4to1_bh mux1(.i(i),.sel(sel),.y(y));

initial
begin
/*	sel = 2'b00; i = 4'b0000;
	#10 i = 4'b0001;
	#10 i = 4'b0010;
	#10 i = 4'b0011;
	#10 i = 4'b0100;
	#10 i = 4'b0101;
	#10 i = 4'b0110;
	#10 i = 4'b0111;
	#10 i = 4'b1000;
	#10 i = 4'b1001;
	#10 i = 4'b1010;
	#10 i = 4'b1011;
	#10 i = 4'b1100;
	#10 i = 4'b1101;
	#10 i = 4'b1110;
	#10 i = 4'b1111;
	#10 sel = 2'b01; i = 4'b0000;
	#10 i = 4'b0001;
	#10 i = 4'b0010;
	#10 i = 4'b0011;
	#10 i = 4'b0100;
	#10 i = 4'b0101;
	#10 i = 4'b0110;
	#10 i = 4'b0111;
	#10 i = 4'b1000;
	#10 i = 4'b1001;
	#10 i = 4'b1010;
	#10 i = 4'b1011;
	#10 i = 4'b1100;
	#10 i = 4'b1101;
	#10 i = 4'b1110;
	#10 i = 4'b1111;
	#10 sel = 2'b10; i = 4'b0000;
	#10 i = 4'b0001;
	#10 i = 4'b0010;
	#10 i = 4'b0011;
	#10 i = 4'b0100;
	#10 i = 4'b0101;
	#10 i = 4'b0110;
	#10 i = 4'b0111;
	#10 i = 4'b1000;
	#10 i = 4'b1001;
	#10 i = 4'b1010;
	#10 i = 4'b1011;
	#10 i = 4'b1100;
	#10 i = 4'b1101;
	#10 i = 4'b1110;
	#10 i = 4'b1111;
	#10 sel = 2'b11; i = 4'b0000;
	#10 i = 4'b0001;
	#10 i = 4'b0010;
	#10 i = 4'b0011;
	#10 i = 4'b0100;
	#10 i = 4'b0101;
	#10 i = 4'b0110;
	#10 i = 4'b0111;
	#10 i = 4'b1000;
	#10 i = 4'b1001;
	#10 i = 4'b1010;
	#10 i = 4'b1011;
	#10 i = 4'b1100;
	#10 i = 4'b1101;
	#10 i = 4'b1110;
	#10 i = 4'b1111; */
	{sel,i} = 6'd0;
	repeat(63)
	#50 {sel,i} = {sel,i} + 1'b1;
end

initial
	$monitor($time," i = %b, sel = %b, y = %b",i,sel,y);

endmodule 