module ha
(input a,b,
 output s,c);

assign s = a^b,
	c = a&b;

endmodule 
