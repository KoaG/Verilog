module test
(input [25:0]i,
output out);

and a1(out,i[25],i[24],i[23],i[22],i[21],i[20],i[19],i[18],i[17],i[16],i[15],i[14],i[13],i[12],i[11],i[10],i[9],i[8],i[7],i[6],i[5],i[4],i[3],i[2],i[1],i[0]);

endmodule 